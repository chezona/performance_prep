`ifndef MEMORY_SYSTOLIC_ARRAY_IF
`define MEMORY_SYSTOLIC_ARRAY_IF

`endif 